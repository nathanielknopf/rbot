// basically need an internal variable that tracks what block of moves to spit out
// can have a memory module that stores a shit ton of strings of moves
// some dumb nerd shit

module spin_all(input send_setup_moves, clock, 
                output reg [n:0] moves);
endmodule